* SPICE3 file created from INVERTOR_TEST_0.ext - technology: sky130A

X0 INV_1445845_0_0_1692204508_0/m1_312_1400# INV_1445845_0_0_1692204508_0/li_405_571# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.294 pd=2.38 as=0.557 ps=4.73 w=2.1 l=0.15
X1 VSUBS INV_1445845_0_0_1692204508_0/li_405_571# INV_1445845_0_0_1692204508_0/m1_312_1400# VSUBS sky130_fd_pr__nfet_01v8 ad=0.557 pd=4.73 as=0.294 ps=2.38 w=2.1 l=0.15
X2 INV_1445845_0_0_1692204508_0/m1_312_1400# INV_1445845_0_0_1692204508_0/li_405_571# INV_1445845_0_0_1692204508_0/PMOS_S_19745913_X1_Y1_1692204509_1692204508_0/w_0_0# INV_1445845_0_0_1692204508_0/PMOS_S_19745913_X1_Y1_1692204509_1692204508_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.38 as=0.557 ps=4.73 w=2.1 l=0.15
X3 INV_1445845_0_0_1692204508_0/PMOS_S_19745913_X1_Y1_1692204509_1692204508_0/w_0_0# INV_1445845_0_0_1692204508_0/li_405_571# INV_1445845_0_0_1692204508_0/m1_312_1400# INV_1445845_0_0_1692204508_0/PMOS_S_19745913_X1_Y1_1692204509_1692204508_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0.557 pd=4.73 as=0.294 ps=2.38 w=2.1 l=0.15
C0 INV_1445845_0_0_1692204508_0/m1_312_1400# INV_1445845_0_0_1692204508_0/li_405_571# 0.241f
C1 INV_1445845_0_0_1692204508_0/li_405_571# INV_1445845_0_0_1692204508_0/PMOS_S_19745913_X1_Y1_1692204509_1692204508_0/w_0_0# 0.89f
C2 INV_1445845_0_0_1692204508_0/m1_312_1400# INV_1445845_0_0_1692204508_0/PMOS_S_19745913_X1_Y1_1692204509_1692204508_0/w_0_0# 0.788f
C3 INV_1445845_0_0_1692204508_0/m1_312_1400# VSUBS 0.898f **FLOATING
C4 INV_1445845_0_0_1692204508_0/li_405_571# VSUBS 1.53f **FLOATING
C5 INV_1445845_0_0_1692204508_0/PMOS_S_19745913_X1_Y1_1692204509_1692204508_0/w_0_0# VSUBS 3.02f **FLOATING
